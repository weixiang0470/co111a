`include "../02/Add16.v"

module main;
reg[15:0] a,b,ans;
wire[15:0] out;
reg[8*1:1] check;

Add16 g0(a,b,out);

//|        a         |        b         |       out        |
//| 0000000000000000 | 0000000000000000 | 0000000000000000 |
//| 0000000000000000 | 1111111111111111 | 1111111111111111 |
//| 1111111111111111 | 1111111111111111 | 1111111111111110 |
//| 1010101010101010 | 0101010101010101 | 1111111111111111 |
//| 0011110011000011 | 0000111111110000 | 0100110010110011 |
//| 0001001000110100 | 1001100001110110 | 1010101010101010 |

initial begin
    $display("\n -------------------------------------------------------------------------");
    $display("|  Time  |         a        |         b         |     Add16Out    | check |");
    $display("|-----------------------------------------------------------------|-------|");
    a=16'b0000000000000000;
    b=16'b0000000000000000;
    ans=16'b0000000000000000;
end
initial #11 begin
    a=16'b0000000000000000;
    b=16'b1111111111111111;
    ans=16'b1111111111111111;
end
initial #21 begin
    a=16'b1111111111111111;
    b=16'b1111111111111111;
    ans=16'b1111111111111110;
end
initial #31 begin
    a=16'b1010101010101010;
    b=16'b0101010101010101;
    ans=16'b1111111111111111;
end
initial #41 begin
    a=16'b0011110011000011;
    b=16'b0000111111110000;
    ans=16'b0100110010110011;
end
initial #51 begin
    a=16'b0001001000110100;
    b=16'b1001100001110110;
    ans=16'b1010101010101010;
end
always #10 begin
    if(out[15:0] == ans[15:0]) check = "v";
    else check="x";
    $display("|%4dns  | %b | %b | %b |   %s   |",$stime,a,b,out,check);
    $display("|-----------------------------------------------------------------|-------|");
end
initial #61 $finish;

endmodule