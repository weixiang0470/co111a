`include "ALU.v"

module main;
reg[15:0] x,y;
reg zx,nx,zy,ny,f,no;
wire[15:0] out;
wire zr,ng;
reg[15:0] Aout;
reg Azr,Ang;
reg[2:0] check;
reg[8*3:1] check2;

ALU g0(x,y,zx,nx,zy,ny,f,no,out,zr,ng);

initial begin
    $display("\n ------------------------------------------------------------------------------------------------|------- ");
    $display("|  Time |        x         |        y         |zx |nx |zy |ny | f |no |       out        |zr |ng | check |");
    $display("|------------------------------------------------------------------------------------------------|-------|");
    x=16'b0000000000000000;y=16'b1111111111111111;
    zx=1;nx=0;zy=1;ny=0;f=1;no=0;
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #11 begin
    zx=1;nx=1;zy=1;ny=1;f=1;no=1;   
    Aout=16'b0000000000000001;Azr=0;Ang=0;
end
initial #21 begin
    zx=1;nx=1;zy=1;ny=0;f=1;no=0;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #31 begin
    zx=0;nx=0;zy=1;ny=1;f=0;no=0;   
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #41 begin
    zx=1;nx=1;zy=0;ny=0;f=0;no=0;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #51 begin
    zx=0;nx=0;zy=1;ny=1;f=0;no=1;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #61 begin
    zx=1;nx=1;zy=0;ny=0;f=0;no=1;   
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #71 begin
    zx=0;nx=0;zy=1;ny=1;f=1;no=1;   
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #81 begin
    zx=1;nx=1;zy=0;ny=0;f=1;no=1;   
    Aout=16'b0000000000000001;Azr=0;Ang=0;
end
initial #91 begin
    zx=0;nx=1;zy=1;ny=1;f=1;no=1;   
    Aout=16'b0000000000000001;Azr=0;Ang=0;
end
initial #101 begin
    zx=1;nx=1;zy=0;ny=1;f=1;no=1;   
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #111 begin
    zx=0;nx=0;zy=1;ny=1;f=1;no=0;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #121 begin
    zx=1;nx=1;zy=0;ny=0;f=1;no=0;   
    Aout=16'b1111111111111110;Azr=0;Ang=1;
end
initial #131 begin
    zx=0;nx=0;zy=0;ny=0;f=1;no=0;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #141 begin
    zx=0;nx=1;zy=0;ny=0;f=1;no=1;   
    Aout=16'b0000000000000001;Azr=0;Ang=0;
end
initial #151 begin
    zx=0;nx=0;zy=0;ny=1;f=1;no=1;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #161 begin
    zx=0;nx=0;zy=0;ny=0;f=0;no=0;   
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #171 begin
    zx=0;nx=1;zy=0;ny=1;f=0;no=1;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #181 begin
    x=16'b0000000000010001;y=16'b0000000000000011;
    zx=1;nx=0;zy=1;ny=0;f=1;no=0;   
    Aout=16'b0000000000000000;Azr=1;Ang=0;
end
initial #191 begin
    zx=1;nx=1;zy=1;ny=1;f=1;no=1;   
    Aout=16'b0000000000000001;Azr=0;Ang=0;
end
initial #201 begin
    zx=1;nx=1;zy=1;ny=0;f=1;no=0;   
    Aout=16'b1111111111111111;Azr=0;Ang=1;
end
initial #211 begin
    zx=0;nx=0;zy=1;ny=1;f=0;no=0;   
    Aout=16'b0000000000010001;Azr=0;Ang=0;
end
initial #221 begin
    zx=1;nx=1;zy=0;ny=0;f=0;no=0;   
    Aout=16'b0000000000000011;Azr=0;Ang=0;
end
initial #231 begin
    zx=0;nx=0;zy=1;ny=1;f=0;no=1;   
    Aout=16'b1111111111101110;Azr=0;Ang=1;
end
initial #241 begin
    zx=1;nx=1;zy=0;ny=0;f=0;no=1;   
    Aout=16'b1111111111111100;Azr=0;Ang=1;
end
initial #251 begin
    zx=0;nx=0;zy=1;ny=1;f=1;no=1;   
    Aout=16'b1111111111101111;Azr=0;Ang=1;
end
initial #261 begin
    zx=1;nx=1;zy=0;ny=0;f=1;no=1;   
    Aout=16'b1111111111111101;Azr=0;Ang=1;
end
initial #271 begin
    zx=0;nx=1;zy=1;ny=1;f=1;no=1;   
    Aout=16'b0000000000010010;Azr=0;Ang=0;
end
initial #281 begin
    zx=1;nx=1;zy=0;ny=1;f=1;no=1;   
    Aout=16'b0000000000000100;Azr=0;Ang=0;
end
initial #291 begin
    zx=0;nx=0;zy=1;ny=1;f=1;no=0;   
    Aout=16'b0000000000010000;Azr=0;Ang=0;
end
initial #301 begin
    zx=1;nx=1;zy=0;ny=0;f=1;no=0;   
    Aout=16'b0000000000000010;Azr=0;Ang=0;
end
initial #311 begin
    zx=0;nx=0;zy=0;ny=0;f=1;no=0;   
    Aout=16'b0000000000010100;Azr=0;Ang=0;
end
initial #321 begin
    zx=0;nx=1;zy=0;ny=0;f=1;no=1;   
    Aout=16'b0000000000001110;Azr=0;Ang=0;
end
initial #331 begin
    zx=0;nx=0;zy=0;ny=1;f=1;no=1;   
    Aout=16'b1111111111110010;Azr=0;Ang=1;
end
initial #341 begin
    zx=0;nx=0;zy=0;ny=0;f=0;no=0;   
    Aout=16'b0000000000000001;Azr=0;Ang=0;
end
initial #351 begin
    zx=0;nx=1;zy=0;ny=1;f=0;no=1;   
    Aout=16'b0000000000010011;Azr=0;Ang=0;
end

initial #361 begin
//1110110000010000
//110000
    x=16'hx;
    y=16'd10;
    zx=1;nx=1;zy=0;ny=0;f=0;no=0;  
    Aout=16'b0000000000001010;Azr=0;Ang=0;
end
always #10 begin
    if(out==Aout)check=4;
    else check=0;
    if(zr==Azr)check=check+2;
    if(ng == Ang)check = check +1;
    if(check==0)check2="xxx";
    if(check==1)check2="xxv";
    if(check==2)check2="xvx";
    if(check==3)check2="xvv";
    if(check==4)check2="vxx";
    if(check==5)check2="vxv";
    if(check==6)check2="vvx";
    if(check==7)check2="vvv";
    $display("|%4dns | %b | %b | %d | %d | %d | %d | %d | %d | %b | %d | %d | %4s  |",$stime,x,y,zx,nx,zy,ny,f,no,out,zr,ng,check2);
    $display("|------------------------------------------------------------------------------------------------|-------|");
end

initial #371 $finish;

endmodule
//---------------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------------------
//|        x         |        y         |zx |nx |zy |ny | f |no |       out        |zr |ng |
//| 0000000000000000 | 1111111111111111 | 1 | 0 | 1 | 0 | 1 | 0 | 0000000000000000 | 1 | 0 | 0ns
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 1 | 1 | 1 | 1 | 0000000000000001 | 0 | 0 | 11ns  
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 1 | 0 | 1 | 0 | 1111111111111111 | 0 | 1 | 21ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 1 | 1 | 0 | 0 | 0000000000000000 | 1 | 0 | 31ns
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 0 | 0 | 0 | 0 | 1111111111111111 | 0 | 1 | 41ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 1 | 1 | 0 | 1 | 1111111111111111 | 0 | 1 | 51ns
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 0 | 0 | 0 | 1 | 0000000000000000 | 1 | 0 | 61ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 1 | 1 | 1 | 1 | 0000000000000000 | 1 | 0 | 71ns
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 0 | 0 | 1 | 1 | 0000000000000001 | 0 | 0 | 81ns
//| 0000000000000000 | 1111111111111111 | 0 | 1 | 1 | 1 | 1 | 1 | 0000000000000001 | 0 | 0 | 91ns
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 0 | 1 | 1 | 1 | 0000000000000000 | 1 | 0 | 101ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 1 | 1 | 1 | 0 | 1111111111111111 | 0 | 1 | 111ns
//| 0000000000000000 | 1111111111111111 | 1 | 1 | 0 | 0 | 1 | 0 | 1111111111111110 | 0 | 1 | 121ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 0 | 0 | 1 | 0 | 1111111111111111 | 0 | 1 | 131ns
//| 0000000000000000 | 1111111111111111 | 0 | 1 | 0 | 0 | 1 | 1 | 0000000000000001 | 0 | 0 | 141ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 0 | 1 | 1 | 1 | 1111111111111111 | 0 | 1 | 151ns
//| 0000000000000000 | 1111111111111111 | 0 | 0 | 0 | 0 | 0 | 0 | 0000000000000000 | 1 | 0 | 161ns
//| 0000000000000000 | 1111111111111111 | 0 | 1 | 0 | 1 | 0 | 1 | 1111111111111111 | 0 | 1 | 171ns
//| 0000000000010001 | 0000000000000011 | 1 | 0 | 1 | 0 | 1 | 0 | 0000000000000000 | 1 | 0 | 181ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 1 | 1 | 1 | 1 | 0000000000000001 | 0 | 0 | 191ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 1 | 0 | 1 | 0 | 1111111111111111 | 0 | 1 | 201ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 1 | 1 | 0 | 0 | 0000000000010001 | 0 | 0 | 211ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 0 | 0 | 0 | 0 | 0000000000000011 | 0 | 0 | 221ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 1 | 1 | 0 | 1 | 1111111111101110 | 0 | 1 | 231ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 0 | 0 | 0 | 1 | 1111111111111100 | 0 | 1 | 241ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 1 | 1 | 1 | 1 | 1111111111101111 | 0 | 1 | 251ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 0 | 0 | 1 | 1 | 1111111111111101 | 0 | 1 | 261ns
//| 0000000000010001 | 0000000000000011 | 0 | 1 | 1 | 1 | 1 | 1 | 0000000000010010 | 0 | 0 | 271ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 0 | 1 | 1 | 1 | 0000000000000100 | 0 | 0 | 281ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 1 | 1 | 1 | 0 | 0000000000010000 | 0 | 0 | 291ns
//| 0000000000010001 | 0000000000000011 | 1 | 1 | 0 | 0 | 1 | 0 | 0000000000000010 | 0 | 0 | 301ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 0 | 0 | 1 | 0 | 0000000000010100 | 0 | 0 | 311ns
//| 0000000000010001 | 0000000000000011 | 0 | 1 | 0 | 0 | 1 | 1 | 0000000000001110 | 0 | 0 | 321ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 0 | 1 | 1 | 1 | 1111111111110010 | 0 | 1 | 331ns
//| 0000000000010001 | 0000000000000011 | 0 | 0 | 0 | 0 | 0 | 0 | 0000000000000001 | 0 | 0 | 341ns
//| 0000000000010001 | 0000000000000011 | 0 | 1 | 0 | 1 | 0 | 1 | 0000000000010011 | 0 | 0 | 351ns
