`include "And16.v"

module main;
reg[15:0] a,b,ans;
wire[15:0] out;

And16 g1(a,b,out);

//|        a         |        b         |       out        |
//| 0000000000000000 | 0000000000000000 | 0000000000000000 |
//| 0000000000000000 | 1111111111111111 | 0000000000000000 |
//| 1111111111111111 | 1111111111111111 | 1111111111111111 |
//| 1010101010101010 | 0101010101010101 | 0000000000000000 |
//| 0011110011000011 | 0000111111110000 | 0000110011000000 |
//| 0001001000110100 | 1001100001110110 | 0001000000110100 |

initial begin
    $display("  Time |        a         |        b         |      And16       |       Ans        |");
    $display("------------------------------------------------------------------------------------");
    $monitor("%4dns | %b | %b | %b | %b |",$stime,a,b,out,ans);
    a=16'b0000000000000000;
    b=16'b0000000000000000;
    ans=16'b0000000000000000;
end

initial #25 begin
    a=16'b0000000000000000;
    b=16'b1111111111111111;
    ans=16'b0000000000000000;
end

initial #50 begin
    a=16'b1111111111111111;
    b=16'b1111111111111111;
    ans=16'b1111111111111111;
end

initial #75 begin
    a=16'b1010101010101010;
    b=16'b0101010101010101;
    ans=16'b0000000000000000;
end

initial #100 begin
    a=16'b0011110011000011;
    b=16'b0000111111110000;
    ans=16'b0000110011000000;
end

initial #125 begin
    a=16'b0001001000110100;
    b=16'b1001100001110110;
    ans=16'b0001000000110100;
end

initial #126 begin
    $display("------------------------------------------------------------------------------------");
end

initial #126 $finish;
endmodule