`include "Mux8Way16.v"

module main;
reg[15:0] d7,d6,d5,d4,d3,d2,d1,d0,ans;
reg[2:0] sel;
wire[15:0] out;
reg[8*1:1] check;

    Mux8Way16 g0(d7,d6,d5,d4,d3,d2,d1,d0,sel,out);

//|        a         |        b         |        c         |        d         |        e         |        f         |        g         |        h         |  sel  |       out        |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  000  | 0001001000110100 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  001  | 0010001101000101 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  010  | 0011010001010110 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  011  | 0100010101100111 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  100  | 0101011001111000 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  101  | 0110011110001001 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  110  | 0111100010011010 |
//| 0001001000110100 | 0010001101000101 | 0011010001010110 | 0100010101100111 | 0101011001111000 | 0110011110001001 | 0111100010011010 | 1000100110101011 |  111  | 1000100110101011 |

initial begin
    d0=16'b0001001000110100;
    d1=16'b0010001101000101;
    d2=16'b0011010001010110;
    d3=16'b0100010101100111;
    d4=16'b0101011001111000;
    d5=16'b0110011110001001;
    d6=16'b0111100010011010;
    d7=16'b1000100110101011;
    $display("\nd0=%b\nd1=%b\nd2=%b\nd3=%b\nd4=%b\nd5=%b\nd6=%b\nd7=%b\n",d0,d1,d2,d3,d4,d5,d6,d7);
    $display(" ----------------------------------------- ");
    $display("|  Time  | sel |     Mux8Way16    | check |");
    $display("|---------------------------------|-------|");
    sel=3'b000;
    ans=16'b0001001000110100;
end
initial #11 begin
    ans=16'b0010001101000101;
end
initial #21 begin
    ans=16'b0011010001010110;
end
initial #31 begin
    ans=16'b0100010101100111;
end
initial #41 begin
    ans=16'b0101011001111000;
end
initial #51 begin
    ans=16'b0110011110001001;
end
initial #61 begin
    ans=16'b0111100010011010;
end
initial #71 begin
    ans=16'b1000100110101011;
end
always #10 begin
    if(out == ans) check="v";
    else check="x";
    $display("|%4dns  | %b | %b | %3s   |",$stime,sel,out,check);
    sel=sel+1;
end
initial #81 begin
    $display(" ----------------------------------------- ");
    #1 $finish;
end

endmodule